LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

package array_machine is
	type logic_array is array (3 downto 0, 4 downto 0) of std_logic;
end array_machine;

package body array_machine is

end array_machine; 